--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   21:26:54 11/09/2016
-- Design Name:   
-- Module Name:   C:/Users/CBAS/Desktop/UTP/Laboratorio de electronica/EJERCICIOS/XILINX PROYECTOS 20152 NOVIEMBRE 07/Procesador4/tb_psr.vhd
-- Project Name:  Procesador4
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: PSR
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY tb_psr IS
END tb_psr;
 
ARCHITECTURE behavior OF tb_psr IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT PSR
    PORT(
         CLK : IN  std_logic;
         Reset : IN  std_logic;
         NZVC : IN  std_logic_vector(3 downto 0);
         Carry : OUT  std_logic;
         NCwp : IN  std_logic;
         Cwp : IN  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal CLK : std_logic := '0';
   signal Reset : std_logic := '0';
   signal NZVC : std_logic_vector(3 downto 0) := (others => '0');
   signal NCwp : std_logic := '0';
   signal Cwp : std_logic := '0';

 	--Outputs
   signal Carry : std_logic;

   -- Clock period definitions
   constant CLK_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: PSR PORT MAP (
          CLK => CLK,
          Reset => Reset,
          NZVC => NZVC,
          Carry => Carry,
          NCwp => NCwp,
          Cwp => Cwp
        );

   -- Clock process definitions
   CLK_process :process
   begin
		CLK <= '0';
		wait for CLK_period/2;
		CLK <= '1';
		wait for CLK_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
  begin		
       Reset <='1';
		NZVC <="0010";
		wait for 50 ns;
		Reset<='0';
		NZVC<="1010";
		wait for 50 ns;
		NZVC<="1110";
		wait for 50 ns;
      NZVC<="0101";

      wait;
   end process;

END;
