--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   21:22:56 11/09/2016
-- Design Name:   
-- Module Name:   C:/Users/CBAS/Desktop/UTP/Laboratorio de electronica/EJERCICIOS/XILINX PROYECTOS 20152 NOVIEMBRE 07/Procesador4/tb_UC.vhd
-- Project Name:  Procesador4
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: UC
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY tb_UC IS
END tb_UC;
 
ARCHITECTURE behavior OF tb_UC IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT UC
    PORT(
         op : IN  std_logic_vector(1 downto 0);
         op3 : IN  std_logic_vector(5 downto 0);
         OutUC : OUT  std_logic_vector(5 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal op : std_logic_vector(1 downto 0) := (others => '0');
   signal op3 : std_logic_vector(5 downto 0) := (others => '0');

 	--Outputs
   signal OutUC : std_logic_vector(5 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
  
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: UC PORT MAP (
          op => op,
          op3 => op3,
          OutUC => OutUC
        );


 

   -- Stimulus process
   stim_proc: process
    begin	

      op <= "10";
		op3<="000000";
		wait for 20 ns;
		op3<="010000";
		wait for 20 ns;
		op3<="011000";
		wait for 20 ns;
		op3<="001000";
		wait for 20 ns;
		op3<="000100";
		wait for 20 ns;
		op3<="010100";
		wait for 20 ns;
		op3<="001100";
		wait for 20 ns;
		op3<="011100";
		wait for 20 ns;
		op3<="000001";
		wait for 20 ns;
		op3<="000101";
		wait for 20 ns;
		op3<="010101";
		wait for 20 ns;
		op3<="010001";
		wait for 20 ns;
		op3<="000010";
		wait for 20 ns;
		op3<="000110";
		wait for 20 ns;
		op3<="010010";
		wait for 20 ns;
		op3<="010110";
		wait for 20 ns;
		op3<="000011";
		wait for 20 ns;
		op3<="000111";
		wait for 20 ns;
		op3<="010011";
		wait for 20 ns;
		op3<="010111";
wait for 20 ns;	
     
   end process;


END;
