----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    22:46:23 10/17/2016 
-- Design Name: 
-- Module Name:    Multiplexor - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Multiplexor is
    Port ( i : in  STD_LOGIC;
           Out_SEU : in  STD_LOGIC_VECTOR (31 downto 0);
           Crs2 : in  STD_LOGIC_VECTOR (31 downto 0);
           Out_MUX : out  STD_LOGIC_VECTOR (31 downto 0));
end Multiplexor;

architecture arq_MUX of Multiplexor is

begin
 process (i,Out_SEU,Crs2)
      begin 
		 if (i='0') then 
		      Out_MUX<=Crs2;
		else
		      if (i='1')then
				     Out_MUX<=Out_SEU;		
            end if;
		end if;
end process	;	

end arq_MUX;

